//======================================================================================
// hdc_top.v - Top-Level Wrapper for HDC Image Classification System
//======================================================================================
//
// DESCRIPTION:
//   Top-level wrapper module providing a clean interface for integrating the HDC
//   classifier into larger FPGA/ASIC systems. This module wraps hdc_classifier.v
//   and provides standardized I/O naming conventions suitable for system integration.
//
// PURPOSE:
//   - System integration wrapper for VIAS (Versatile Image Analysis System)
//   - Provides standardized signal naming (pix_in, conf_in, etc.)
//   - Maps between top-level conventions and hdc_classifier interface
//   - Reserved interfaces for future features (scan chain, status registers)
//
// KEY FEATURES:
//   - Direct pass-through to hdc_classifier core
//   - All parameters exposed for flexibility
//   - SystemVerilog 'logic' type for cleaner syntax
//   - Reserved scan chain interface (DFT placeholder)
//   - Status output for system monitoring
//
// USAGE IN SYSTEM:
//   1. Instantiate in top-level FPGA/ASIC design
//   2. Connect clk_in to system clock
//   3. Load configuration via conf_valid_in/conf_in serial interface
//   4. Stream images via pix_in with write_enable pulse
//   5. Read predictions from predicted_class when valid_out asserts
//
// VERIFIED CONFIGURATION (Manufacturing Dataset):
//   - ROW_SZ = 32, HEIGHT_SZ = 32, ADC_BIT_WIDTH = 16
//   - NUM_CLASSES = 2, HDC_HV_DIM = 5000
//   - Achieves 98% accuracy on manufacturing inspection data
//
// AUTHORS:
//   Created by: George Michelogiannakis (mihelog@lbl.gov)
//   Developed with assistance from AI tools (Claude and Gemini)
//   Lawrence Berkeley National Laboratory
//   Created: 2025-09-02
//
//======================================================================================

module hdc_top #(
    //==================================================================================
    // IMAGE PARAMETERS
    //==================================================================================
    parameter ROW_SZ = 32,                           // Image width in pixels (X-axis)
    parameter HEIGHT_SZ = 32,                        // Image height in pixels (Y-axis)
    parameter ADC_BIT_WIDTH = 8,                     // Bits per pixel (8 or 16-bit)

    //==================================================================================
    // CLASSIFICATION PARAMETERS
    //==================================================================================
    parameter NUM_CLASSES = 2,                       // Number of output classes (2-100)
    parameter HDC_HV_DIM = 5000,                     // Hypervector dimension (1000-10000)
    parameter HDC_CONF_WIDTH = 4,                    // Confidence bits (4 = 0-15 range)
    parameter CONFIDENCE_LUT_SIZE = 5000,            // Confidence LUT entries (match HV_DIM)
    parameter ENABLE_ONLINE_LEARNING = 1,            // Enable online learning (0=off, 1=on)
                                                     // This parameter enables OL logic synthesis
                                                     // Actual OL enable controlled by config bit
    parameter CLASS_WIDTH = $clog2(NUM_CLASSES),     // Bits to encode class ID (auto-calculated)

    //==================================================================================
    // CNN WEIGHT PARAMETERS (Must match Python training)
    //==================================================================================
    parameter CONV1_WEIGHT_WIDTH = 12,               // Conv1 weight bit width (8-16 bits)
    parameter CONV2_WEIGHT_WIDTH = 10,               // Conv2 weight bit width (8-16 bits)
    parameter FC_WEIGHT_WIDTH = 8,                   // FC weight bit width (8-bit for 70KB target, 2026-02-04)
    parameter FC_BIAS_WIDTH = 8,                     // FC bias bit width (8-bit for precision, 2026-02-03)
    parameter WEIGHT_WIDTH = 16,                     // General weight width (legacy)

    //==================================================================================
    // QUANTIZATION SCALE PARAMETERS (Generated by Python QAT training)
    // These scales map floating-point weights to fixed-point integers
    //==================================================================================
    parameter real CONV1_WEIGHT_SCALE = 512.0,       // Conv1 weight quantization scale
    parameter real CONV1_BIAS_SCALE = 512.0,         // Conv1 bias quantization scale
    parameter real CONV2_WEIGHT_SCALE = 128.0,       // Conv2 weight quantization scale
    parameter real CONV2_BIAS_SCALE = 128.0,         // Conv2 bias quantization scale
    parameter real FC_WEIGHT_SCALE = 32.0,           // FC weight quantization scale
    parameter real FC_BIAS_SCALE = 64.0,             // FC bias quantization scale

    //==================================================================================
    // PARALLELISM PARAMETERS (Performance tuning)
    // Higher values = faster processing, more area
    //==================================================================================
    parameter PARALLEL_PROJ = 20,                    // Projection dims/cycle (1-100)
    parameter PARALLEL_CONV1 = 8,                    // Conv1 parallel channels (1, 2, 4, 8)
    parameter PARALLEL_CONV2 = 4,                    // Conv2 parallel channels (1, 2, 4, 8, 16)

    //==================================================================================
    // HDC PARAMETERS
    //==================================================================================
    parameter FC_OUT_SIZE = 64,                      // FC layer output size (64 or 128, default: 64)
    parameter HDC_PROJ_WEIGHT_WIDTH = 4,             // Projection weight bits (1, 3, 4, 8)
    parameter ENCODING_LEVELS = 4,                   // Encoding levels (3=ternary, 4=quaternary)
    parameter USE_PER_FEATURE_THRESHOLDS = 1,        // 1=per-feature thresholds, 0=global thresholds
    parameter USE_LFSR_PROJECTION = 0,               // 1=on-the-fly LFSR projection, 0=stored matrix
    parameter LFSR_MASTER_SEED = 32'd42              // Master seed for LFSR (seed[i] = MASTER_SEED + i + 1)
) (
    //==================================================================================
    // CLOCK AND RESET (Synchronous interface)
    //==================================================================================
    input logic reset_b,                             // Active-low asynchronous reset
    input logic clk_in,                              // System clock (100-500 MHz typical)

    //==================================================================================
    // SCAN CHAIN INTERFACE (Reserved for Design-for-Test)
    // Currently unused - placeholder for future DFT features
    //==================================================================================
    input logic scan_en,                             // Scan chain enable (DFT mode)
    input logic scan_clk,                            // Scan chain clock
    input logic scan_in,                             // Scan chain data input
    output logic scan_out,                           // Scan chain data output

    //==================================================================================
    // CONFIGURATION INTERFACE (Serial bitstream loading)
    //==================================================================================
    input logic conf_valid_in,                       // Configuration write enable
                                                     // Assert to load config bits serially
    input logic conf_in,                             // Configuration data bit
                                                     // Serial stream of weights & hypervectors

    //==================================================================================
    // IMAGE INPUT INTERFACE
    //==================================================================================
    input write_enable,                              // Image valid signal (start classification)
                                                     // Pulse high to process pix_in
    input logic [ROW_SZ*ROW_SZ*ADC_BIT_WIDTH-1:0] pix_in,
                                                     // Flattened input image (row-major order)
                                                     // For 32×32×16: [16383:0] = 1024 pixels

    //==================================================================================
    // CLASSIFICATION OUTPUT INTERFACE
    //==================================================================================
    output logic [CLASS_WIDTH-1:0] predicted_class,  // Predicted class ID
                                                     // Valid when valid_out asserts
    output logic [HDC_CONF_WIDTH-1:0] confidence,    // Confidence score (0-15)
                                                     // Higher = more confident
    output logic valid_out,                          // Output valid flag
                                                     // Asserts when classification complete

    //==================================================================================
    // STATUS INTERFACE
    //==================================================================================
    output logic loading_complete,                   // Config loading complete flag
                                                     // Asserts when ready to classify
    output logic ready,                              // Ready for new image flag
                                                     // Asserts when pipeline idle
    output logic [7:0] status                        // General status output
                                                     // Currently fixed at 0xE (example)
);

//======================================================================================
// INTERNAL PARAMETERS
//======================================================================================
localparam shortint LENGTH = 64;                     // Scan chain length (reserved for DFT)

//======================================================================================
// MODULE INSTANTIATION - HDC Classifier Core
//======================================================================================
// Instantiate the main HDC classifier module
// All top-level parameters are passed through to the core
// Signal mappings:
//   - conf_valid_in → write_enable (config loading)
//   - write_enable → valid (image classification trigger)
//   - clk_in → clk (main system clock)
//======================================================================================
hdc_classifier #(
    .IMG_WIDTH(ROW_SZ),
    .IMG_HEIGHT(HEIGHT_SZ),
    .PIXEL_WIDTH(ADC_BIT_WIDTH),
    .NUM_CLASSES(NUM_CLASSES),
    .FC_OUT_SIZE(FC_OUT_SIZE),
    .HDC_HV_DIM(HDC_HV_DIM),
    .HDC_CONF_WIDTH(HDC_CONF_WIDTH),
    .CONFIDENCE_LUT_SIZE(CONFIDENCE_LUT_SIZE),
    .CONV1_WEIGHT_WIDTH(CONV1_WEIGHT_WIDTH),
    .CONV2_WEIGHT_WIDTH(CONV2_WEIGHT_WIDTH),
    .FC_WEIGHT_WIDTH(FC_WEIGHT_WIDTH),
    .FC_BIAS_WIDTH(FC_BIAS_WIDTH),
    .WEIGHT_WIDTH(WEIGHT_WIDTH),
    .CONV1_WEIGHT_SCALE(CONV1_WEIGHT_SCALE),
    .CONV1_BIAS_SCALE(CONV1_BIAS_SCALE),
    .CONV2_WEIGHT_SCALE(CONV2_WEIGHT_SCALE),
    .CONV2_BIAS_SCALE(CONV2_BIAS_SCALE),
    .FC_WEIGHT_SCALE(FC_WEIGHT_SCALE),
    .FC_BIAS_SCALE(FC_BIAS_SCALE),
    .ENABLE_ONLINE_LEARNING(ENABLE_ONLINE_LEARNING),
    .PARALLEL_PROJ(PARALLEL_PROJ),
    .PARALLEL_CONV1(PARALLEL_CONV1),
    .PARALLEL_CONV2(PARALLEL_CONV2),
    .HDC_PROJ_WEIGHT_WIDTH(HDC_PROJ_WEIGHT_WIDTH),
    .ENCODING_LEVELS(ENCODING_LEVELS),
    .USE_PER_FEATURE_THRESHOLDS(USE_PER_FEATURE_THRESHOLDS),
    .USE_LFSR_PROJECTION(USE_LFSR_PROJECTION),
    .LFSR_MASTER_SEED(LFSR_MASTER_SEED)
) hdc_classifier_instance (
    //==================================================================================
    // Clock and Reset
    //==================================================================================
    .clk(clk_in),                                    // Map clk_in → clk
    .reset_b(reset_b),                               // Direct connection

    //==================================================================================
    // Image Classification Interface
    //==================================================================================
    .valid(write_enable),                            // Map write_enable → valid
                                                     // Signals start of classification
    .image_data(pix_in),                             // Direct image input connection

    //==================================================================================
    // Configuration Loading Interface
    //==================================================================================
    .write_enable(conf_valid_in),                    // Map conf_valid_in → write_enable
                                                     // Controls serial config loading
    .data_in(conf_in),                               // Serial configuration bitstream

    //==================================================================================
    // Classification Output Interface
    //==================================================================================
    .predicted_class(predicted_class),               // Direct connection
    .confidence(confidence),                         // Direct connection
    .valid_out(valid_out),                           // Direct connection
    .loading_complete(loading_complete),             // Direct connection
    .ready(ready)                                    // Direct connection
);


//======================================================================================
// INTERNAL SIGNALS
//======================================================================================
logic [LENGTH-1:0] scan_data;                        // Scan chain data buffer (unused)

//======================================================================================
// SCAN CHAIN INSTANTIATION (Currently Commented Out)
//======================================================================================
// Reserved for future Design-for-Test (DFT) implementation
// Uncomment when scan chain testing is needed
//
//scan_chain #(
//    .LENGTH (LENGTH)
//) scan_chain (
//    .reset_b  (reset_b),
//    .scan_en  (scan_en),
//    .scan_clk (scan_clk),
//    .scan_in  (scan_in),
//    .scan_out (scan_out),
//    .scan_data (scan_data)
//);

//======================================================================================
// STATUS OUTPUT
//======================================================================================
// Example status output - currently fixed value
// Can be extended for system monitoring:
//   - Bit 0: Loading complete
//   - Bit 1: Classification active
//   - Bit 2: Online learning active
//   - Bit 3: Error flag
//   - Bits 7-4: Reserved
assign status = 8'hE;                                // Fixed status (0000_1110)


endmodule //hdc_top
